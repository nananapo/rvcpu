`ifndef PKG_CONF_H
`define PKG_CONF_H

package conf;
parameter FREQUENCY_MHz = 27;
parameter UART_BAUDRATE = 115200;
endpackage

`endif