module GlobalHistory2bit #(
    parameter WIDTH_PC = 20,
    parameter WIDTH_HIST = 20
)(
    input wire          clk,
    input wire [31:0]   pc,         // 予測したいアドレス
    output wire [31:0]  next_pc,    // pcから予測された次のアドレス
    input wire IUpdatePredictionIO updateio
);

localparam SIZE_PC = 2 ** WIDTH_PC;
localparam SIZE_HIST = 2 ** WIDTH_HIST;

localparam DEFAULT_COUNTER_VALUE = 2'b0;
localparam DEFAULT_HISTORY_VALUE = {WIDTH_HIST{1'b0}};

logic [1:0]  counters [SIZE_HIST-1:0]; // hist -> counter
logic [31:0] targets [SIZE_PC-1:0]; // pc -> target

initial begin
    for (int i = 0; i < SIZE_HIST; i++)
        counters[i] = DEFAULT_COUNTER_VALUE;
end

logic [WIDTH_HIST-1:0] hist = DEFAULT_HISTORY_VALUE; 

wire [WIDTH_PC-1:0] pci   = pc[WIDTH_PC+2-1:2];
wire [WIDTH_PC-1:0] u_pci = updateio.pc[WIDTH_PC+2-1:2];

// TODO フェッチした時のhistが欲しいが、持ってこれない
wire [1:0] count    = counters[hist];
wire [1:0] u_count  = counters[hist]; // ここ

wire [31:0] target_untaken = pc + 4;
wire [31:0] target_taken   = targets[pci];
assign next_pc = count[1] == 1'b1 ? target_taken : target_untaken;

always @(posedge clk) begin
    if (updateio.valid) begin
        hist <= {hist[WIDTH_HIST-2:0], updateio.taken};

        if (updateio.taken) begin
            targets[u_pci] <= updateio.target;
        end

        if (!(u_count == 2'b11 && updateio.taken) && 
            !(u_count == 2'b00 && !updateio.taken)) begin
            if (updateio.taken)
                counters[hist] <= u_count + 2'b1;
            else
                counters[hist] <= u_count - 2'b1;
        end
    end
end

/*
`ifdef PRINT_DEBUGINFO
always @(posedge clk) begin
    $display("data,fetchstage.glbh2.pc,h,%b", pc);
    $display("data,fetchstage.glbh2.pci,h,%b", pci);
    $display("data,fetchstage.glbh2.hist,b,%b", hist);
    $display("data,fetchstage.glbh2.count,b,%b", count);
    $display("data,fetchstage.glbh2.next_pc,h,%b", next_pc);
end
`endif 
*/

endmodule