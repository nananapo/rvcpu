module CSRStage(
	input wire clk
);



endmodule